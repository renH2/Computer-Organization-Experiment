`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:17:10 08/15/2020 
// Design Name: 
// Module Name:    Mul32 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Mul32(
	input clk,
	input [31:0]A,B,
	input Ctrl,//�����з��Ż����޷��ų˳�
	output reg [63:0]Mul_Out
    );
	 reg [61:0]mul_out;

	 reg [30:0]C,D;	 
	 always@(*)begin
	 if(A[31]==1'b1)
		C<=(~A[30:0])+1;
	 else
		C<=A[30:0];
	 if(B[31]==1'b1)
		D<=(~B[30:0])+1;
	 else
		D<=B[30:0];
	 case(Ctrl)
	 1'b0:begin
    Mul_Out<={32'b00000000000000000000000000000000, {32{B[0]}}&A       }+{31'b0000000000000000000000000000000, {32{B[1]}}&A, 1'b0  }+{30'b000000000000000000000000000000, {32{B[2]}}&A, 2'b00  }+{29'b00000000000000000000000000000, {32{B[3]}}&A, 3'b000  }
				+{28'b0000000000000000000000000000, {32{B[4]}}&A, 4'b0000  }+{27'b000000000000000000000000000, {32{B[5]}}&A, 5'b00000  }+{26'b00000000000000000000000000, {32{B[6]}}&A, 6'b000000  }+{25'b0000000000000000000000000, {32{B[7]}}&A, 7'b0000000  }
				+{24'b000000000000000000000000, {32{B[8]}}&A, 8'b00000000  }+{23'b00000000000000000000000, {32{B[9]}}&A, 9'b000000000  }+{22'b0000000000000000000000, {32{B[10]}}&A, 10'b0000000000}+{21'b000000000000000000000, {32{B[11]}}&A, 11'b00000000000}
				+{20'b00000000000000000000, {32{B[12]}}&A, 12'b000000000000}+{19'b0000000000000000000, {32{B[13]}}&A, 13'b0000000000000}+{18'b000000000000000000, {32{B[14]}}&A, 14'b00000000000000}+{17'b00000000000000000, {32{B[15]}}&A, 15'b000000000000000}
				+{16'b0000000000000000, {32{B[16]}}&A, 16'b0000000000000000}+{15'b000000000000000, {32{B[17]}}&A, 17'b00000000000000000}+{14'b00000000000000, {32{B[18]}}&A, 18'b000000000000000000}+{13'b0000000000000, {32{B[19]}}&A, 19'b0000000000000000000}
				+{12'b000000000000, {32{B[20]}}&A, 20'b00000000000000000000}+{11'b00000000000, {32{B[21]}}&A, 21'b000000000000000000000}+{10'b0000000000, {32{B[22]}}&A, 22'b0000000000000000000000}+{9'b000000000, {32{B[23]}}&A, 23'b00000000000000000000000 }
				+{ 8'b00000000, {32{B[24]}}&A, 24'b000000000000000000000000}+{7'b0000000, {32{B[25]}}&A, 25'b0000000000000000000000000 }+{6'b000000, {32{B[26]}}&A, 26'b00000000000000000000000000 }+{5'b00000, {32{B[27]}}&A, 27'b000000000000000000000000000 }
				+{ 4'b0000, {32{B[28]}}&A, 28'b0000000000000000000000000000}+{3'b000, {32{B[29]}}&A, 29'b00000000000000000000000000000 }+{2'b00, {32{B[30]}}&A, 30'b000000000000000000000000000000 }+{1'b0, {32{B[31]}}&A, 31'b0000000000000000000000000000000 };
			end
	1'b1:begin
	/*mul_out<={31'b0000000000000000000000000000000, {31{B[0]}}&A[30:0] }+{30'b000000000000000000000000000000, {31{B[1]}}&A[30:0] ,1'b0}+{29'b00000000000000000000000000000, {31{B[2]}}&A[30:0] ,2'b00}+{28'b0000000000000000000000000000, {31{B[3]}}&A[30:0] ,3'b000}
			  +{27'b000000000000000000000000000, {31{B[4]}}&A[30:0] ,4'b0000}+{26'b00000000000000000000000000, {31{B[5]}}&A[30:0] ,5'b00000}+{25'b0000000000000000000000000, {31{B[6]}}&A[30:0] ,6'b000000}+{24'b000000000000000000000000, {31{B[7]}}&A[30:0] ,7'b0000000}
			  +{23'b00000000000000000000000, {31{B[8]}}&A[30:0] ,8'b00000000}+{22'b0000000000000000000000, {31{B[9]}}&A[30:0] ,9'b000000000}+{21'b000000000000000000000, {31{B[10]}}&A[30:0] ,10'b0000000000}+{20'b00000000000000000000, {31{B[11]}}&A[30:0] ,11'b00000000000}
			  +{19'b0000000000000000000, {31{B[12]}}&A[30:0] ,12'b000000000000}+{18'b000000000000000000, {31{B[13]}}&A[30:0] ,13'b0000000000000}+{17'b00000000000000000, {31{B[14]}}&A[30:0] ,14'b00000000000000}+{16'b0000000000000000, {31{B[15]}}&A[30:0] ,15'b000000000000000}
			  +{15'b000000000000000, {31{B[16]}}&A[30:0] ,16'b0000000000000000}+{14'b00000000000000, {31{B[17]}}&A[30:0] ,17'b00000000000000000}+{13'b0000000000000, {31{B[18]}}&A[30:0] ,18'b000000000000000000}+{12'b000000000000, {31{B[19]}}&A[30:0] ,19'b0000000000000000000}
			  +{11'b00000000000, {31{B[20]}}&A[30:0] ,20'b00000000000000000000}+{10'b0000000000, {31{B[21]}}&A[30:0] ,21'b000000000000000000000}+{9'b000000000, {31{B[22]}}&A[30:0] ,22'b0000000000000000000000}+{8'b00000000, {31{B[23]}}&A[30:0] ,23'b00000000000000000000000}
			  +{7'b0000000, {31{B[24]}}&A[30:0] ,24'b000000000000000000000000}+{6'b000000, {31{B[25]}}&A[30:0] ,25'b0000000000000000000000000}+{5'b00000, {31{B[26]}}&A[30:0] ,26'b00000000000000000000000000}+{4'b0000, {31{B[27]}}&A[30:0] ,27'b000000000000000000000000000}
			  +{3'b000, {31{B[28]}}&A[30:0] ,28'b0000000000000000000000000000}+{2'b00, {31{B[29]}}&A[30:0] ,29'b00000000000000000000000000000}+{1'b0, {31{B[30]}}&A[30:0] ,30'b000000000000000000000000000000};
*/	
	mul_out<={31'b0000000000000000000000000000000,{31{D[0]}}&C[30:0]}+{30'b000000000000000000000000000000,{31{D[1]}}&C[30:0],1'b0}+{29'b00000000000000000000000000000,{31{D[2]}}&C[30:0],2'b00}+{28'b0000000000000000000000000000,{31{D[3]}}&C[30:0],3'b000}
			  +{27'b000000000000000000000000000,{31{D[4]}}&C[30:0],4'b0000}+{26'b00000000000000000000000000,{31{D[5]}}&C[30:0],5'b00000}+{25'b0000000000000000000000000,{31{D[6]}}&C[30:0],6'b000000}+{24'b000000000000000000000000,{31{D[7]}}&C[30:0],7'b0000000}
			  +{23'b00000000000000000000000,{31{D[8]}}&C[30:0],8'b00000000}+{22'b0000000000000000000000,{31{D[9]}}&C[30:0],9'b000000000}+{21'b000000000000000000000,{31{D[10]}}&C[30:0],10'b0000000000}+{20'b00000000000000000000,{31{D[11]}}&C[30:0],11'b00000000000}
			  +{19'b0000000000000000000,{31{D[12]}}&C[30:0],12'b000000000000}+{18'b000000000000000000,{31{D[13]}}&C[30:0],13'b0000000000000}+{17'b00000000000000000,{31{D[14]}}&C[30:0],14'b00000000000000}+{16'b0000000000000000,{31{D[15]}}&C[30:0],15'b000000000000000}
			  +{15'b000000000000000,{31{D[16]}}&C[30:0],16'b0000000000000000}+{14'b00000000000000,{31{D[17]}}&C[30:0],17'b00000000000000000}+{13'b0000000000000,{31{D[18]}}&C[30:0],18'b000000000000000000}+{12'b000000000000,{31{D[19]}}&C[30:0],19'b0000000000000000000}
			  +{11'b00000000000,{31{D[20]}}&C[30:0],20'b00000000000000000000}+{10'b0000000000,{31{D[21]}}&C[30:0],21'b000000000000000000000}+{9'b000000000,{31{D[22]}}&C[30:0],22'b0000000000000000000000}+{8'b00000000,{31{D[23]}}&C[30:0],23'b00000000000000000000000}
			  +{7'b0000000,{31{D[24]}}&C[30:0],24'b000000000000000000000000}+{6'b000000,{31{D[25]}}&C[30:0],25'b0000000000000000000000000}+{5'b00000,{31{D[26]}}&C[30:0],26'b00000000000000000000000000}+{4'b0000,{31{D[27]}}&C[30:0],27'b000000000000000000000000000}
			  +{3'b000,{31{D[28]}}&C[30:0],28'b0000000000000000000000000000}+{2'b00,{31{D[29]}}&C[30:0],29'b00000000000000000000000000000}+{1'b0,{31{D[30]}}&C[30:0],30'b000000000000000000000000000000};
	Mul_Out<={A[31]^B[31],1'b0,mul_out}; 
			  end
	endcase
	end
endmodule
